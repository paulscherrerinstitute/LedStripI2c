library ieee;

use ieee.std_logic_1164.all;

package MpcI2cSequencerPkg is 

  -- if CTRL is '1' and last is '0'  then a restart is generated
  -- if CTRL and LAST are both set then a STOP is generated

  constant MPCI2C_CTRL_C : natural := 8;
  constant MPCI2C_LAST_C : natural := 9;
  constant MPCI2C_RDNW_C : natural := 0;

  -- prepend any of these to a data byte;
  -- If the bus is not currently held, the first item (even if SEQ_NORM) generates a start condition
  -- and therefore the associated data must be a bus address + R/W bit.
  constant SEQ_NORM        : std_logic_vector(1 downto 0) := "00"; -- data byte to send
  constant SEQ_RSRT        : std_logic_vector(1 downto 0) := "01"; -- restart; data is bus address + R/W
  constant SEQ_LAST        : std_logic_vector(1 downto 0) := "10"; -- last byte to send; no STOP
  constant SEQ_STOP        : std_logic_vector(1 downto 0) := "11"; -- last byte to send; STOP

  subtype  MpcI2cSequenceDataType is std_logic_vector(MPCI2C_LAST_C downto 0);

  type     MpcI2cSequenceArray    is array(natural range<>) of MpcI2cSequenceDataType;

  -- An I2C Sequencer program is a sequence of 10-bit values:
  --
  --  LAST_BIT, CTRL_BIT, DATA_BITS(7 downto 0)
  --
  -- 1. A START condition is generated by
  --     - the first element in a sequence
  --     - an element which has the CTRL_BIT set and LAST_BIT clear
  --       (RESTART).
  --
  --   DATA_BITS(7 downto 1) define the target i2c address
  --   and DATA_BITS(0) the direction of the subsequent data
  --   transfers ('1' -> READ, '0' -> WRITE).
  --
  -- 2. In WRITE mode (sequence elements following a START
  --    or RESTART element) DATA_BITS(7 downto 0) are sent over I2C.
  --
  -- 3. In READ mode the sequence element following a START or
  --    RESTART element defines the number of bytes to read from
  --    the target.
  --     num_bytes : DATA_BITS(7 downto 0) + 1
  --    If LAST_BIT is clear and CTRL_BIT is set then the last
  --    byte is NOT acknowledged by the master. This is useful
  --    if more than 256 bytes need to be read, e.g., 
  --
  --      "01" & "1010000" & "1" -- RESTART a READ from address 0x50
  --      "01" & x"ff"           -- read 256 bytes (no final NACK)
  --      "00" & x"00"           -- read one more byte, send NAK
  --
  -- If the LAST_BIT is asserted then this flags an element as the
  -- last element of a sequence, i.e., no more subsequent elments
  -- are fetched and executed.
  -- If the CTRL_BIT is asserted together with LAST then a STOP condition
  -- is generated. If CTRL_BIT is clear then the bus is kept.
  --
  -- Example:
  --
  --     "00" & "1010000" & "0" -- START (first element) a WRITE to address 0x50
  --     "00" & x"00"           -- WRITE 0x00
  --     "01" & "1010000" & "1" -- RESTART a READ from address 0x50
  --     "10" & x"04"           -- READ 5 bytes, generate NAK, terminate program
  --                            -- but keep the bus
  --     "01" & "1010000" & "0" -- RESTART write to address 0x50 (new program)
  --     "11" & x"00"           -- WRITE 0, generate STOP and terminate program
  --
  --     Note that the above memory contents define two separate programs
  --     that need to be passed to the controller separately:
  --
  --     signal memPtr      : natural   := 0;
  --     signal memPtrValid : std_logic := '1';
  --
  --     if ( rising_edge(clk) ) then
  --       if ( (memPtrReady = '1') and (memPtrValid = '1') ) then
  --         if ( memPtr = 0 ) then
  --            -- second program
  --            memPtr <= 4; -- offset of 2nd program
  --         else
  --            memPtrValid <= '0';
  --         end if;
  --       end if;
  --     end if;
  -- 

end package MpcI2cSequencerPkg;
